

library IEEE;
use IEEE.STD_LOGIC_1164.all;

package Pack is
type memArray64 is array(0 to 63) of std_logic_vector(31 downto 0);
type memArray8 is array(0 to 7) of std_logic_vector(31 downto 0);


end Pack;

package body Pack is
 
end Pack;
