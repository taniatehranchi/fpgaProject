library IEEE;
use IEEE.STD_LOGIC_1164.all;

package matrix is
type matrix64 is array(0 to 63) of std_logic_vector(31 downto 0);
type matrix8 is array(0 to 7) of std_logic_vector(31 downto 0);


end matrix;

package body matrix is
 
end matrix;
